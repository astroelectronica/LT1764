.title KiCad schematic
.include "C:/AE/LT1764/_models/C3216X5R2A105K160AA_s.mod"
.include "C:/AE/LT1764/_models/CGA5L3X5R1H106K160AB_s.mod"
.include "C:/AE/LT1764/_models/LT1764.lib"
V1 /VIN 0 {VSOURCE}
XU2 /VOUT /ADJ 0 /VIN /VIN LT1764MD
XU1 /VIN 0 C3216X5R2A105K160AA_s
R2 /VOUT /ADJ {RADJU}
R3 /ADJ 0 {RADJB}
I1 /VOUT 0 {ILOAD}
XU3 /VOUT 0 CGA5L3X5R1H106K160AB_s
.end
